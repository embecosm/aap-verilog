module Clock (CLOCK_50, clock);

	output clock;
	input CLOCK_50;
	
	wire clock = CLOCK_50;
	
endmodule
